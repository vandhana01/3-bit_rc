magic
tech sky130A
magscale 1 2
timestamp 1700904678
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 2128 98808 97424
<< metal2 >>
rect 61198 99200 61254 100000
rect 18 0 74 800
rect 77942 0 77998 800
<< obsm2 >>
rect 20 99144 61142 99362
rect 61310 99144 98422 99362
rect 20 856 98422 99144
rect 130 800 77886 856
rect 78054 800 98422 856
<< metal3 >>
rect 0 82288 800 82408
rect 99200 58488 100000 58608
<< obsm3 >>
rect 800 82488 99200 97409
rect 880 82208 99200 82488
rect 800 58688 99200 82208
rect 800 58408 99120 58688
rect 800 2143 99200 58408
<< metal4 >>
rect 1944 2128 2264 97424
rect 2604 2128 2924 97424
rect 6944 2128 7264 97424
rect 7604 2128 7924 97424
rect 11944 2128 12264 97424
rect 12604 2128 12924 97424
rect 16944 2128 17264 97424
rect 17604 2128 17924 97424
rect 21944 2128 22264 97424
rect 22604 2128 22924 97424
rect 26944 2128 27264 97424
rect 27604 2128 27924 97424
rect 31944 2128 32264 97424
rect 32604 2128 32924 97424
rect 36944 2128 37264 97424
rect 37604 2128 37924 97424
rect 41944 2128 42264 97424
rect 42604 2128 42924 97424
rect 46944 2128 47264 97424
rect 47604 2128 47924 97424
rect 51944 2128 52264 97424
rect 52604 2128 52924 97424
rect 56944 2128 57264 97424
rect 57604 2128 57924 97424
rect 61944 2128 62264 97424
rect 62604 2128 62924 97424
rect 66944 2128 67264 97424
rect 67604 2128 67924 97424
rect 71944 2128 72264 97424
rect 72604 2128 72924 97424
rect 76944 2128 77264 97424
rect 77604 2128 77924 97424
rect 81944 2128 82264 97424
rect 82604 2128 82924 97424
rect 86944 2128 87264 97424
rect 87604 2128 87924 97424
rect 91944 2128 92264 97424
rect 92604 2128 92924 97424
rect 96944 2128 97264 97424
rect 97604 2128 97924 97424
<< metal5 >>
rect 1056 93676 98856 93996
rect 1056 93016 98856 93336
rect 1056 88676 98856 88996
rect 1056 88016 98856 88336
rect 1056 83676 98856 83996
rect 1056 83016 98856 83336
rect 1056 78676 98856 78996
rect 1056 78016 98856 78336
rect 1056 73676 98856 73996
rect 1056 73016 98856 73336
rect 1056 68676 98856 68996
rect 1056 68016 98856 68336
rect 1056 63676 98856 63996
rect 1056 63016 98856 63336
rect 1056 58676 98856 58996
rect 1056 58016 98856 58336
rect 1056 53676 98856 53996
rect 1056 53016 98856 53336
rect 1056 48676 98856 48996
rect 1056 48016 98856 48336
rect 1056 43676 98856 43996
rect 1056 43016 98856 43336
rect 1056 38676 98856 38996
rect 1056 38016 98856 38336
rect 1056 33676 98856 33996
rect 1056 33016 98856 33336
rect 1056 28676 98856 28996
rect 1056 28016 98856 28336
rect 1056 23676 98856 23996
rect 1056 23016 98856 23336
rect 1056 18676 98856 18996
rect 1056 18016 98856 18336
rect 1056 13676 98856 13996
rect 1056 13016 98856 13336
rect 1056 8676 98856 8996
rect 1056 8016 98856 8336
rect 1056 3676 98856 3996
rect 1056 3016 98856 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42604 2128 42924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47604 2128 47924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 52604 2128 52924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57604 2128 57924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 62604 2128 62924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67604 2128 67924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 72604 2128 72924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 77604 2128 77924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 82604 2128 82924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 87604 2128 87924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 92604 2128 92924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97604 2128 97924 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 98856 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 98856 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 98856 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 98856 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 98856 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 98856 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 98856 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 38676 98856 38996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43676 98856 43996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 48676 98856 48996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 53676 98856 53996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 58676 98856 58996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 63676 98856 63996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 68676 98856 68996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 73676 98856 73996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 78676 98856 78996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 83676 98856 83996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 88676 98856 88996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 93676 98856 93996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41944 2128 42264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46944 2128 47264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 51944 2128 52264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 56944 2128 57264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 61944 2128 62264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 66944 2128 67264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 71944 2128 72264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 76944 2128 77264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 81944 2128 82264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 86944 2128 87264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 91944 2128 92264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96944 2128 97264 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 98856 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 98856 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 98856 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 98856 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 98856 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 98856 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 98856 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 38016 98856 38336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 43016 98856 43336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 48016 98856 48336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 53016 98856 53336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 58016 98856 58336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 63016 98856 63336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 68016 98856 68336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 73016 98856 73336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 78016 98856 78336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 83016 98856 83336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 88016 98856 88336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 93016 98856 93336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 82288 800 82408 6 clk
port 3 nsew signal input
rlabel metal2 s 18 0 74 800 6 count[0]
port 4 nsew signal output
rlabel metal3 s 99200 58488 100000 58608 6 count[1]
port 5 nsew signal output
rlabel metal2 s 61198 99200 61254 100000 6 count[2]
port 6 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 ori
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5473970
string GDS_FILE /home/vandhana/3-bit_rc/openlane/pes_3bit_rc/runs/23_11_25_14_58/results/signoff/pes_3bit_rc.magic.gds
string GDS_START 102176
<< end >>

