VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pes_3bit_rc
  CLASS BLOCK ;
  FOREIGN pes_3bit_rc ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.020 10.640 114.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 10.640 139.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.020 10.640 164.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 10.640 189.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.020 10.640 214.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 10.640 239.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.020 10.640 264.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.020 10.640 289.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 313.020 10.640 314.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 10.640 339.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 363.020 10.640 364.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 10.640 389.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.020 10.640 414.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.020 10.640 439.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 463.020 10.640 464.620 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.020 10.640 489.620 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 494.280 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 494.280 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 494.280 69.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 93.380 494.280 94.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 118.380 494.280 119.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 143.380 494.280 144.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 168.380 494.280 169.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 193.380 494.280 194.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 218.380 494.280 219.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 243.380 494.280 244.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 268.380 494.280 269.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 293.380 494.280 294.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 318.380 494.280 319.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 343.380 494.280 344.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 368.380 494.280 369.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 393.380 494.280 394.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 418.380 494.280 419.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 443.380 494.280 444.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 468.380 494.280 469.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.720 10.640 111.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 10.640 136.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 10.640 161.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 10.640 186.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.720 10.640 211.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 10.640 236.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.720 10.640 261.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.720 10.640 286.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.720 10.640 311.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 10.640 336.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.720 10.640 361.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 10.640 386.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 409.720 10.640 411.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.720 10.640 436.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.720 10.640 461.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.720 10.640 486.320 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 494.280 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 494.280 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 494.280 66.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 90.080 494.280 91.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 115.080 494.280 116.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 140.080 494.280 141.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 165.080 494.280 166.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 190.080 494.280 191.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 215.080 494.280 216.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 240.080 494.280 241.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 265.080 494.280 266.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 290.080 494.280 291.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 315.080 494.280 316.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 340.080 494.280 341.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 365.080 494.280 366.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 390.080 494.280 391.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 415.080 494.280 416.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 440.080 494.280 441.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 465.080 494.280 466.680 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END count[0]
  PIN count[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END count[1]
  PIN count[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 305.990 496.000 306.270 500.000 ;
    END
  END count[2]
  PIN ori
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END ori
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 0.100 495.720 305.710 496.810 ;
        RECT 306.550 495.720 492.110 496.810 ;
        RECT 0.100 4.280 492.110 495.720 ;
        RECT 0.650 4.000 389.430 4.280 ;
        RECT 390.270 4.000 492.110 4.280 ;
      LAYER met3 ;
        RECT 4.000 412.440 496.000 487.045 ;
        RECT 4.400 411.040 496.000 412.440 ;
        RECT 4.000 293.440 496.000 411.040 ;
        RECT 4.000 292.040 495.600 293.440 ;
        RECT 4.000 10.715 496.000 292.040 ;
  END
END pes_3bit_rc
END LIBRARY

